`timescale 1ns/100ps
/*
Title         :  CIC Filter
Project       :  tt06

Filename      :  CIC.v
Author        :  Madeline Crowley
Created       :  04/06/2024 16:44:39
Last Modified :  04/06/2024 16:46:37
Copyright (c) :  Madeline (Liam) Crowley

INPUTS        :
OUTPUTS       :
PARAMETERS    :

Description   : Cascaded integrator-comb variable filter

Mod History   : 04/06/2024 16:44:39 : created
*/

module CIC (
    // Ports
);



endmodule: CIC
