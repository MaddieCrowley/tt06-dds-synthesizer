`timescale 1ns/100ps
/*
Title         :  tb_Filter
Project       :  tt06

Filename      :  tb_Filter.v
Author        :  Madeline Crowley
Created       :  03/02/2024 18:57:58
Last Modified :  03/02/2024 18:58:30
Copyright (c) :  Madeline (Liam) Crowley

INPUTS        : 
OUTPUTS       : 
PARAMETERS    : 

Description   : Testbench for the filter module

Mod History   : 03/02/2024 18:57:58 : created
*/

